
module c432 ( N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, 
        N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, 
        N89, N92, N95, N99, N102, N105, N108, N112, N115, N223, N329, N370, 
        N421, N430, N431, N432 );
  input N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47,
         N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92,
         N95, N99, N102, N105, N108, N112, N115;
  output N223, N329, N370, N421, N430, N431, N432;
  wire   N203, N309, N360, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209;
  assign N223 = N203;
  assign N329 = N309;
  assign N370 = N360;

  HDOAI21DL U100 ( .A1(n117), .A2(n118), .B(n119), .Z(N432) );
  HDAOI21D1 U101 ( .A1(n120), .A2(n121), .B(n122), .Z(n118) );
  HDOAI21DL U102 ( .A1(n123), .A2(n124), .B(n125), .Z(n122) );
  HDINVBD1 U103 ( .A(n126), .Z(n123) );
  HDINVBD1 U104 ( .A(n127), .Z(n117) );
  HDNAN3D1 U105 ( .A1(n119), .A2(n127), .A3(n128), .Z(N431) );
  HDNAN3D1 U106 ( .A1(n126), .A2(n129), .A3(n125), .Z(n128) );
  HDOA32DL U107 ( .A1(N430), .A2(n120), .A3(n130), .B1(n131), .B2(n132), .Z(
        N421) );
  HDAO22DL U108 ( .A1(N309), .A2(N8), .B1(N360), .B2(N14), .Z(n132) );
  HDOAI21DL U109 ( .A1(n133), .A2(n134), .B(n135), .Z(n130) );
  HDINVBD1 U110 ( .A(n129), .Z(n135) );
  HDNAN2D1 U111 ( .A1(n124), .A2(n121), .Z(n129) );
  HDOAI222DL U112 ( .A1(n136), .A2(n137), .B1(n138), .B2(n139), .C1(n140), 
        .C2(n141), .Z(n121) );
  HDNOR2D1 U113 ( .A1(N203), .A2(n142), .Z(n140) );
  HDINVBD1 U114 ( .A(N92), .Z(n139) );
  HDINVBD1 U115 ( .A(N86), .Z(n137) );
  HDAO211DL U116 ( .A1(N360), .A2(N79), .B(n143), .C(n144), .Z(n124) );
  HDAO21DL U117 ( .A1(N73), .A2(N309), .B(n145), .Z(n144) );
  HDOAI21DL U118 ( .A1(n136), .A2(n146), .B(N108), .Z(n134) );
  HDOAI21DL U119 ( .A1(n138), .A2(n147), .B(n148), .Z(n133) );
  HDINVBD1 U120 ( .A(N115), .Z(n147) );
  HDAOI222D1 U121 ( .A1(n149), .A2(n150), .B1(N309), .B2(N99), .C1(N360), .C2(
        N105), .Z(n120) );
  HDNAN2D1 U122 ( .A1(n151), .A2(N95), .Z(n149) );
  HDNAN4D1 U123 ( .A1(n125), .A2(n126), .A3(n119), .A4(n127), .Z(N430) );
  HDOAI211DL U124 ( .A1(n138), .A2(n152), .B(n153), .C(n154), .Z(n127) );
  HDAOI21D1 U125 ( .A1(N24), .A2(N203), .B(n155), .Z(n154) );
  HDINVBD1 U126 ( .A(N40), .Z(n152) );
  HDOAI211DL U127 ( .A1(n138), .A2(n156), .B(n157), .C(n158), .Z(n119) );
  HDAOI21D1 U128 ( .A1(N21), .A2(N309), .B(n159), .Z(n158) );
  HDOAI211DL U129 ( .A1(n138), .A2(n160), .B(n161), .C(n162), .Z(n126) );
  HDAOI21D1 U130 ( .A1(N60), .A2(N309), .B(n163), .Z(n162) );
  HDINVBD1 U131 ( .A(N66), .Z(n160) );
  HDINVBD1 U132 ( .A(N360), .Z(n138) );
  HDAO211DL U133 ( .A1(N360), .A2(N53), .B(n164), .C(n165), .Z(n125) );
  HDAO21DL U134 ( .A1(N47), .A2(N309), .B(n166), .Z(n165) );
  HDNAN4D1 U135 ( .A1(n167), .A2(n168), .A3(n169), .A4(n170), .Z(N360) );
  HDNOR3DL U136 ( .A1(n171), .A2(n172), .A3(n173), .Z(n170) );
  HDNOR3DL U137 ( .A1(n174), .A2(N53), .A3(n164), .Z(n173) );
  HDOAI21DL U138 ( .A1(n175), .A2(n136), .B(N43), .Z(n174) );
  HDNOR4M1DL U139 ( .A1(n153), .A2(N40), .A3(n176), .A4(n155), .Z(n172) );
  HDNAN2D1 U140 ( .A1(N34), .A2(N309), .Z(n153) );
  HDOAI31DL U141 ( .A1(n177), .A2(N79), .A3(n143), .B(n178), .Z(n171) );
  HDOAI211DL U142 ( .A1(n179), .A2(n151), .B(N56), .C(n180), .Z(n178) );
  HDAOI21D1 U143 ( .A1(N309), .A2(n181), .B(N66), .Z(n180) );
  HDINVBD1 U144 ( .A(N50), .Z(n179) );
  HDOAI21DL U145 ( .A1(n182), .A2(n136), .B(N69), .Z(n177) );
  HDAOI21D1 U146 ( .A1(n183), .A2(n184), .B(n185), .Z(n169) );
  HDOAI33DL U147 ( .A1(n186), .A2(N92), .A3(n187), .B1(n188), .B2(N105), .B3(
        n189), .Z(n185) );
  HDOAI21DL U148 ( .A1(n190), .A2(n136), .B(N95), .Z(n188) );
  HDOAI21DL U149 ( .A1(n191), .A2(n136), .B(N82), .Z(n186) );
  HDAOI21D1 U150 ( .A1(N309), .A2(n192), .B(N115), .Z(n184) );
  HDAOI21D1 U151 ( .A1(N203), .A2(N102), .B(n193), .Z(n183) );
  HDOAI211DL U152 ( .A1(n194), .A2(n151), .B(N4), .C(n195), .Z(n168) );
  HDAOI21D1 U153 ( .A1(N8), .A2(N309), .B(N14), .Z(n195) );
  HDNAN3D1 U154 ( .A1(n157), .A2(n156), .A3(n196), .Z(n167) );
  HDOA21DL U155 ( .A1(n197), .A2(n136), .B(N17), .Z(n196) );
  HDINVBD1 U156 ( .A(N309), .Z(n136) );
  HDINVBD1 U157 ( .A(N27), .Z(n156) );
  HDNAN4D1 U158 ( .A1(n181), .A2(n192), .A3(n198), .A4(n199), .Z(N309) );
  HDNOR3DL U159 ( .A1(n200), .A2(n175), .A3(n197), .Z(n199) );
  HDNOR3M1DL U160 ( .A1(n157), .A2(N21), .A3(n159), .Z(n197) );
  HDNAN2M1D1 U161 ( .A1(n201), .A2(N203), .Z(n157) );
  HDNOR3DL U162 ( .A1(n164), .A2(N47), .A3(n166), .Z(n175) );
  HDNOR2D1 U163 ( .A1(n151), .A2(n202), .Z(n164) );
  HDOAI32DL U164 ( .A1(n155), .A2(N34), .A3(n176), .B1(N8), .B2(n131), .Z(n200) );
  HDOAI21DL U165 ( .A1(n151), .A2(n194), .B(N4), .Z(n131) );
  HDINVBD1 U166 ( .A(N1), .Z(n194) );
  HDAND2D1 U167 ( .A1(N24), .A2(N203), .Z(n176) );
  HDNOR3DL U168 ( .A1(n190), .A2(n182), .A3(n191), .Z(n198) );
  HDNOR3DL U169 ( .A1(n187), .A2(N86), .A3(n142), .Z(n191) );
  HDNOR2D1 U170 ( .A1(n151), .A2(n141), .Z(n187) );
  HDNOR3DL U171 ( .A1(n143), .A2(N73), .A3(n145), .Z(n182) );
  HDNOR2D1 U172 ( .A1(n151), .A2(n203), .Z(n143) );
  HDNOR3DL U173 ( .A1(n189), .A2(N99), .A3(n204), .Z(n190) );
  HDNOR2D1 U174 ( .A1(n151), .A2(n205), .Z(n189) );
  HDINVBD1 U175 ( .A(N203), .Z(n151) );
  HDNAN3D1 U176 ( .A1(n148), .A2(n146), .A3(N108), .Z(n192) );
  HDINVBD1 U177 ( .A(N112), .Z(n146) );
  HDNAN2D1 U178 ( .A1(N102), .A2(N203), .Z(n148) );
  HDNAN3M1DL U179 ( .A1(N60), .A2(n161), .A3(N56), .Z(n181) );
  HDNAN2D1 U180 ( .A1(N50), .A2(N203), .Z(n161) );
  HDNAN4M1DL U181 ( .A1(n141), .A2(n150), .A3(n206), .A4(n207), .Z(N203) );
  HDNOR2D1 U182 ( .A1(n208), .A2(n209), .Z(n207) );
  HDOAI22DL U183 ( .A1(N50), .A2(n163), .B1(N24), .B2(n155), .Z(n209) );
  HDINVBD1 U184 ( .A(N30), .Z(n155) );
  HDINVBD1 U185 ( .A(N56), .Z(n163) );
  HDOAI22M10D1 U186 ( .A1(N4), .A2(N1), .B1(N102), .B2(n193), .Z(n208) );
  HDINVBD1 U187 ( .A(N108), .Z(n193) );
  HDNOR3DL U188 ( .A1(n201), .A2(n203), .A3(n202), .Z(n206) );
  HDNOR2D1 U189 ( .A1(N37), .A2(n166), .Z(n202) );
  HDINVBD1 U190 ( .A(N43), .Z(n166) );
  HDNOR2D1 U191 ( .A1(N63), .A2(n145), .Z(n203) );
  HDINVBD1 U192 ( .A(N69), .Z(n145) );
  HDNOR2D1 U193 ( .A1(N11), .A2(n159), .Z(n201) );
  HDINVBD1 U194 ( .A(N17), .Z(n159) );
  HDINVBD1 U195 ( .A(n205), .Z(n150) );
  HDNOR2D1 U196 ( .A1(N89), .A2(n204), .Z(n205) );
  HDINVBD1 U197 ( .A(N95), .Z(n204) );
  HDNOR2D1 U198 ( .A1(N76), .A2(n142), .Z(n141) );
  HDINVBD1 U199 ( .A(N82), .Z(n142) );
endmodule

