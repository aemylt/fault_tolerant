
module c499 ( N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, 
        N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, 
        N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, 
        N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, 
        N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, 
        N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
  input N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57,
         N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109,
         N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135,
         N136, N137;
  output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734,
         N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745,
         N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
  wire   n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259;

  HDOA33D1 U157 ( .A1(n160), .A2(n185), .A3(n162), .B1(n165), .B2(n186), .B3(
        n157), .Z(n139) );
  HDOA33D1 U158 ( .A1(n177), .A2(n176), .A3(n178), .B1(n167), .B2(n166), .B3(
        n168), .Z(n140) );
  HDEXOR2D1 U159 ( .A1(N125), .A2(n141), .Z(N755) );
  HDNOR2D1 U160 ( .A1(n142), .A2(n143), .Z(n141) );
  HDEXOR2D1 U161 ( .A1(N121), .A2(n144), .Z(N754) );
  HDNOR2D1 U162 ( .A1(n145), .A2(n143), .Z(n144) );
  HDEXOR2D1 U163 ( .A1(N117), .A2(n146), .Z(N753) );
  HDNOR2D1 U164 ( .A1(n147), .A2(n143), .Z(n146) );
  HDEXOR2D1 U165 ( .A1(N113), .A2(n148), .Z(N752) );
  HDNOR2D1 U166 ( .A1(n149), .A2(n143), .Z(n148) );
  HDNAN3D1 U167 ( .A1(n150), .A2(n151), .A3(n152), .Z(n143) );
  HDNOR3DL U168 ( .A1(n153), .A2(n139), .A3(n154), .Z(n152) );
  HDEXNOR2D1 U169 ( .A1(N109), .A2(n155), .Z(N751) );
  HDNAN2D1 U170 ( .A1(n156), .A2(n157), .Z(n155) );
  HDEXOR2D1 U171 ( .A1(n158), .A2(n159), .Z(N750) );
  HDNAN2D1 U172 ( .A1(n156), .A2(n160), .Z(n159) );
  HDEXNOR2D1 U173 ( .A1(N101), .A2(n161), .Z(N749) );
  HDNAN2D1 U174 ( .A1(n156), .A2(n162), .Z(n161) );
  HDEXOR2D1 U175 ( .A1(n163), .A2(n164), .Z(N748) );
  HDNAN2D1 U176 ( .A1(n156), .A2(n165), .Z(n164) );
  HDNOR4M1DL U177 ( .A1(n166), .A2(n167), .A3(n168), .A4(n139), .Z(n156) );
  HDEXNOR2D1 U178 ( .A1(N93), .A2(n169), .Z(N747) );
  HDNAN2D1 U179 ( .A1(n170), .A2(n157), .Z(n169) );
  HDEXOR2D1 U180 ( .A1(n171), .A2(n172), .Z(N746) );
  HDNAN2D1 U181 ( .A1(n170), .A2(n160), .Z(n172) );
  HDEXOR2D1 U182 ( .A1(n173), .A2(n174), .Z(N745) );
  HDNAN2D1 U183 ( .A1(n170), .A2(n162), .Z(n174) );
  HDEXNOR2D1 U184 ( .A1(N81), .A2(n175), .Z(N744) );
  HDNAN2D1 U185 ( .A1(n170), .A2(n165), .Z(n175) );
  HDNOR4M1DL U186 ( .A1(n176), .A2(n177), .A3(n178), .A4(n139), .Z(n170) );
  HDEXOR2D1 U187 ( .A1(N77), .A2(n179), .Z(N743) );
  HDNOR2D1 U188 ( .A1(n142), .A2(n180), .Z(n179) );
  HDEXOR2D1 U189 ( .A1(N73), .A2(n181), .Z(N742) );
  HDNOR2D1 U190 ( .A1(n145), .A2(n180), .Z(n181) );
  HDEXOR2D1 U191 ( .A1(N69), .A2(n182), .Z(N741) );
  HDNOR2D1 U192 ( .A1(n147), .A2(n180), .Z(n182) );
  HDEXOR2D1 U193 ( .A1(N65), .A2(n183), .Z(N740) );
  HDNOR2D1 U194 ( .A1(n149), .A2(n180), .Z(n183) );
  HDNAN3D1 U195 ( .A1(n153), .A2(n154), .A3(n184), .Z(n180) );
  HDNOR3DL U196 ( .A1(n151), .A2(n139), .A3(n150), .Z(n184) );
  HDEXOR2D1 U197 ( .A1(N61), .A2(n187), .Z(N739) );
  HDNOR2D1 U198 ( .A1(n153), .A2(n188), .Z(n187) );
  HDEXOR2D1 U199 ( .A1(N57), .A2(n189), .Z(N738) );
  HDNOR2D1 U200 ( .A1(n151), .A2(n188), .Z(n189) );
  HDEXOR2D1 U201 ( .A1(N53), .A2(n190), .Z(N737) );
  HDNOR2D1 U202 ( .A1(n154), .A2(n188), .Z(n190) );
  HDEXOR2D1 U203 ( .A1(N49), .A2(n191), .Z(N736) );
  HDNOR2D1 U204 ( .A1(n150), .A2(n188), .Z(n191) );
  HDNAN3D1 U205 ( .A1(n149), .A2(n145), .A3(n192), .Z(n188) );
  HDNOR3DL U206 ( .A1(n142), .A2(n140), .A3(n147), .Z(n192) );
  HDEXNOR2D1 U207 ( .A1(N45), .A2(n193), .Z(N735) );
  HDNAN2D1 U208 ( .A1(n194), .A2(n167), .Z(n193) );
  HDEXNOR2D1 U209 ( .A1(N41), .A2(n195), .Z(N734) );
  HDNAN2D1 U210 ( .A1(n194), .A2(n178), .Z(n195) );
  HDEXOR2D1 U211 ( .A1(n196), .A2(n197), .Z(N733) );
  HDNAN2D1 U212 ( .A1(n194), .A2(n177), .Z(n197) );
  HDEXNOR2D1 U213 ( .A1(N33), .A2(n198), .Z(N732) );
  HDNAN2D1 U214 ( .A1(n194), .A2(n168), .Z(n198) );
  HDNOR4M1DL U215 ( .A1(n186), .A2(n165), .A3(n157), .A4(n140), .Z(n194) );
  HDINVBD1 U216 ( .A(n142), .Z(n157) );
  HDINVBD1 U217 ( .A(n149), .Z(n165) );
  HDNOR2D1 U218 ( .A1(n147), .A2(n145), .Z(n186) );
  HDEXOR2D1 U219 ( .A1(n199), .A2(n200), .Z(N731) );
  HDNAN2D1 U220 ( .A1(n201), .A2(n167), .Z(n200) );
  HDEXNOR2D1 U221 ( .A1(N25), .A2(n202), .Z(N730) );
  HDNAN2D1 U222 ( .A1(n201), .A2(n178), .Z(n202) );
  HDEXNOR2D1 U223 ( .A1(N21), .A2(n203), .Z(N729) );
  HDNAN2D1 U224 ( .A1(n201), .A2(n177), .Z(n203) );
  HDEXOR2D1 U225 ( .A1(n204), .A2(n205), .Z(N728) );
  HDNAN2D1 U226 ( .A1(n201), .A2(n168), .Z(n205) );
  HDNOR4M1DL U227 ( .A1(n185), .A2(n160), .A3(n162), .A4(n140), .Z(n201) );
  HDINVBD1 U228 ( .A(n147), .Z(n162) );
  HDINVBD1 U229 ( .A(n145), .Z(n160) );
  HDNOR2D1 U230 ( .A1(n142), .A2(n149), .Z(n185) );
  HDEXOR2D1 U231 ( .A1(N13), .A2(n206), .Z(N727) );
  HDNOR2D1 U232 ( .A1(n153), .A2(n207), .Z(n206) );
  HDEXOR2D1 U233 ( .A1(N9), .A2(n208), .Z(N726) );
  HDNOR2D1 U234 ( .A1(n151), .A2(n207), .Z(n208) );
  HDEXOR2D1 U235 ( .A1(N5), .A2(n209), .Z(N725) );
  HDNOR2D1 U236 ( .A1(n154), .A2(n207), .Z(n209) );
  HDEXOR2D1 U237 ( .A1(N1), .A2(n210), .Z(N724) );
  HDNOR2D1 U238 ( .A1(n150), .A2(n207), .Z(n210) );
  HDNAN3D1 U239 ( .A1(n147), .A2(n142), .A3(n211), .Z(n207) );
  HDNOR3DL U240 ( .A1(n149), .A2(n140), .A3(n145), .Z(n211) );
  HDEXOR3D1 U241 ( .A1(n212), .A2(n213), .A3(n214), .Z(n145) );
  HDEXOR2D1 U242 ( .A1(n215), .A2(n216), .Z(n214) );
  HDNAN2D1 U243 ( .A1(N137), .A2(N135), .Z(n215) );
  HDEXOR3D1 U244 ( .A1(N121), .A2(N105), .A3(n217), .Z(n213) );
  HDEXOR2D1 U245 ( .A1(N89), .A2(N73), .Z(n217) );
  HDINVBD1 U246 ( .A(n150), .Z(n168) );
  HDNOR2D1 U247 ( .A1(n151), .A2(n154), .Z(n166) );
  HDINVBD1 U248 ( .A(n153), .Z(n167) );
  HDINVBD1 U249 ( .A(n151), .Z(n178) );
  HDEXOR3D1 U250 ( .A1(n218), .A2(n219), .A3(n220), .Z(n151) );
  HDEXOR2D1 U251 ( .A1(n221), .A2(n222), .Z(n220) );
  HDNAN2D1 U252 ( .A1(N131), .A2(N137), .Z(n221) );
  HDEXOR3D1 U253 ( .A1(N41), .A2(N25), .A3(n223), .Z(n219) );
  HDEXOR2D1 U254 ( .A1(N9), .A2(N57), .Z(n223) );
  HDNOR2D1 U255 ( .A1(n153), .A2(n150), .Z(n176) );
  HDEXOR3D1 U256 ( .A1(n224), .A2(n225), .A3(n226), .Z(n153) );
  HDEXOR2D1 U257 ( .A1(n227), .A2(n228), .Z(n226) );
  HDNAN2D1 U258 ( .A1(N132), .A2(N137), .Z(n227) );
  HDEXOR3D1 U259 ( .A1(N29), .A2(N13), .A3(n229), .Z(n225) );
  HDEXOR2D1 U260 ( .A1(N61), .A2(N45), .Z(n229) );
  HDINVBD1 U261 ( .A(n154), .Z(n177) );
  HDEXOR3D1 U262 ( .A1(n222), .A2(n230), .A3(n231), .Z(n154) );
  HDEXOR2D1 U263 ( .A1(n232), .A2(n228), .Z(n231) );
  HDEXNOR3D1 U264 ( .A1(N117), .A2(N113), .A3(n233), .Z(n228) );
  HDEXNOR2D1 U265 ( .A1(N121), .A2(N125), .Z(n233) );
  HDNAN2D1 U266 ( .A1(N130), .A2(N137), .Z(n232) );
  HDEXOR3D1 U267 ( .A1(N37), .A2(N21), .A3(n234), .Z(n230) );
  HDEXOR2D1 U268 ( .A1(N53), .A2(N5), .Z(n234) );
  HDEXOR3D1 U269 ( .A1(n158), .A2(N101), .A3(n235), .Z(n222) );
  HDEXOR2D1 U270 ( .A1(N109), .A2(n163), .Z(n235) );
  HDINVBD1 U271 ( .A(N97), .Z(n163) );
  HDINVBD1 U272 ( .A(N105), .Z(n158) );
  HDEXOR3D1 U273 ( .A1(n212), .A2(n236), .A3(n237), .Z(n149) );
  HDEXOR2D1 U274 ( .A1(n238), .A2(n239), .Z(n237) );
  HDNAN2D1 U275 ( .A1(N133), .A2(N137), .Z(n238) );
  HDEXOR3D1 U276 ( .A1(N65), .A2(N113), .A3(n240), .Z(n236) );
  HDEXOR2D1 U277 ( .A1(N97), .A2(N81), .Z(n240) );
  HDEXNOR3D1 U278 ( .A1(N13), .A2(N1), .A3(n241), .Z(n212) );
  HDEXNOR2D1 U279 ( .A1(N5), .A2(N9), .Z(n241) );
  HDEXOR3D1 U280 ( .A1(n239), .A2(n242), .A3(n243), .Z(n142) );
  HDEXOR2D1 U281 ( .A1(n244), .A2(n245), .Z(n243) );
  HDNAN2D1 U282 ( .A1(N136), .A2(N137), .Z(n244) );
  HDEXOR3D1 U283 ( .A1(N125), .A2(N109), .A3(n246), .Z(n242) );
  HDEXOR2D1 U284 ( .A1(N93), .A2(N77), .Z(n246) );
  HDEXOR3D1 U285 ( .A1(N21), .A2(n204), .A3(n247), .Z(n239) );
  HDEXOR2D1 U286 ( .A1(N25), .A2(n199), .Z(n247) );
  HDINVBD1 U287 ( .A(N29), .Z(n199) );
  HDINVBD1 U288 ( .A(N17), .Z(n204) );
  HDEXOR3D1 U289 ( .A1(n216), .A2(n248), .A3(n249), .Z(n147) );
  HDEXOR2D1 U290 ( .A1(n250), .A2(n245), .Z(n249) );
  HDEXNOR3D1 U291 ( .A1(N53), .A2(N49), .A3(n251), .Z(n245) );
  HDEXNOR2D1 U292 ( .A1(N57), .A2(N61), .Z(n251) );
  HDNAN2D1 U293 ( .A1(N134), .A2(N137), .Z(n250) );
  HDEXOR3D1 U294 ( .A1(N117), .A2(N101), .A3(n252), .Z(n248) );
  HDEXOR2D1 U295 ( .A1(N85), .A2(N69), .Z(n252) );
  HDEXOR3D1 U296 ( .A1(n196), .A2(N33), .A3(n253), .Z(n216) );
  HDEXNOR2D1 U297 ( .A1(N41), .A2(N45), .Z(n253) );
  HDINVBD1 U298 ( .A(N37), .Z(n196) );
  HDEXOR3D1 U299 ( .A1(n218), .A2(n254), .A3(n255), .Z(n150) );
  HDEXOR2D1 U300 ( .A1(n256), .A2(n224), .Z(n255) );
  HDEXOR3D1 U301 ( .A1(n173), .A2(N81), .A3(n257), .Z(n224) );
  HDEXOR2D1 U302 ( .A1(n171), .A2(N93), .Z(n257) );
  HDINVBD1 U303 ( .A(N89), .Z(n171) );
  HDINVBD1 U304 ( .A(N85), .Z(n173) );
  HDNAN2D1 U305 ( .A1(N129), .A2(N137), .Z(n256) );
  HDEXOR3D1 U306 ( .A1(N17), .A2(N1), .A3(n258), .Z(n254) );
  HDEXOR2D1 U307 ( .A1(N49), .A2(N33), .Z(n258) );
  HDEXNOR3D1 U308 ( .A1(N69), .A2(N65), .A3(n259), .Z(n218) );
  HDEXNOR2D1 U309 ( .A1(N73), .A2(N77), .Z(n259) );
endmodule

