
module c1355 ( G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, 
        G1329, G1330, G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, 
        G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, G1348, 
        G1349, G1350, G1351, G1352, G1353, G1354, G1355, G14, G15, G16, G17, 
        G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
        G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, 
        G7, G8, G9 );
  input G1, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G2, G20, G21,
         G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34,
         G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9;
  output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333,
         G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343,
         G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353,
         G1354, G1355;
  wire   n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352;

  HDEXNOR2D1 U201 ( .A1(G32), .A2(n211), .Z(G1355) );
  HDNOR2D1 U202 ( .A1(n212), .A2(n213), .Z(n211) );
  HDEXOR2D1 U203 ( .A1(n214), .A2(n215), .Z(G1354) );
  HDNOR2D1 U204 ( .A1(n216), .A2(n213), .Z(n215) );
  HDEXNOR2D1 U205 ( .A1(G30), .A2(n217), .Z(G1353) );
  HDNOR2D1 U206 ( .A1(n218), .A2(n213), .Z(n217) );
  HDEXNOR2D1 U207 ( .A1(G29), .A2(n219), .Z(G1352) );
  HDNOR2D1 U208 ( .A1(n220), .A2(n213), .Z(n219) );
  HDNAN3D1 U209 ( .A1(n221), .A2(n222), .A3(n223), .Z(n213) );
  HDNOR3DL U210 ( .A1(n224), .A2(n225), .A3(n226), .Z(n223) );
  HDEXOR2D1 U211 ( .A1(n227), .A2(G28), .Z(G1351) );
  HDNAN2D1 U212 ( .A1(n228), .A2(n229), .Z(n227) );
  HDEXOR2D1 U213 ( .A1(n230), .A2(G27), .Z(G1350) );
  HDNAN2D1 U214 ( .A1(n228), .A2(n231), .Z(n230) );
  HDEXOR2D1 U215 ( .A1(n232), .A2(G26), .Z(G1349) );
  HDNAN2D1 U216 ( .A1(n228), .A2(n233), .Z(n232) );
  HDEXOR2D1 U217 ( .A1(n234), .A2(G25), .Z(G1348) );
  HDNAN2D1 U218 ( .A1(n228), .A2(n235), .Z(n234) );
  HDNOR4M1DL U219 ( .A1(n236), .A2(n221), .A3(n226), .A4(n225), .Z(n228) );
  HDEXOR2D1 U220 ( .A1(n237), .A2(G24), .Z(G1347) );
  HDNAN2D1 U221 ( .A1(n238), .A2(n229), .Z(n237) );
  HDEXOR2D1 U222 ( .A1(n239), .A2(G23), .Z(G1346) );
  HDNAN2D1 U223 ( .A1(n238), .A2(n231), .Z(n239) );
  HDEXOR2D1 U224 ( .A1(n240), .A2(G22), .Z(G1345) );
  HDNAN2D1 U225 ( .A1(n238), .A2(n233), .Z(n240) );
  HDEXOR2D1 U226 ( .A1(n241), .A2(G21), .Z(G1344) );
  HDNAN2D1 U227 ( .A1(n238), .A2(n235), .Z(n241) );
  HDNOR4M1DL U228 ( .A1(n242), .A2(n222), .A3(n224), .A4(n225), .Z(n238) );
  HDEXNOR2D1 U229 ( .A1(G20), .A2(n243), .Z(G1343) );
  HDNOR2D1 U230 ( .A1(n212), .A2(n244), .Z(n243) );
  HDEXOR2D1 U231 ( .A1(n245), .A2(n246), .Z(G1342) );
  HDNOR2D1 U232 ( .A1(n216), .A2(n244), .Z(n246) );
  HDEXNOR2D1 U233 ( .A1(G18), .A2(n247), .Z(G1341) );
  HDNOR2D1 U234 ( .A1(n218), .A2(n244), .Z(n247) );
  HDEXNOR2D1 U235 ( .A1(G17), .A2(n248), .Z(G1340) );
  HDNOR2D1 U236 ( .A1(n220), .A2(n244), .Z(n248) );
  HDNAN3D1 U237 ( .A1(n224), .A2(n226), .A3(n249), .Z(n244) );
  HDNOR3DL U238 ( .A1(n222), .A2(n225), .A3(n221), .Z(n249) );
  HDOA33D1 U239 ( .A1(n233), .A2(n250), .A3(n231), .B1(n229), .B2(n251), .B3(
        n235), .Z(n225) );
  HDEXNOR2D1 U240 ( .A1(G16), .A2(n252), .Z(G1339) );
  HDNOR2D1 U241 ( .A1(n253), .A2(n254), .Z(n252) );
  HDEXOR2D1 U242 ( .A1(n255), .A2(n256), .Z(G1338) );
  HDNOR2D1 U243 ( .A1(n257), .A2(n254), .Z(n256) );
  HDEXNOR2D1 U244 ( .A1(G14), .A2(n258), .Z(G1337) );
  HDNOR2D1 U245 ( .A1(n259), .A2(n254), .Z(n258) );
  HDEXOR2D1 U246 ( .A1(n260), .A2(n261), .Z(G1336) );
  HDNOR2D1 U247 ( .A1(n262), .A2(n254), .Z(n261) );
  HDNAN3D1 U248 ( .A1(n233), .A2(n229), .A3(n263), .Z(n254) );
  HDNOR3DL U249 ( .A1(n235), .A2(n264), .A3(n231), .Z(n263) );
  HDEXOR2D1 U250 ( .A1(n265), .A2(G12), .Z(G1335) );
  HDNAN2D1 U251 ( .A1(n266), .A2(n221), .Z(n265) );
  HDEXOR2D1 U252 ( .A1(n267), .A2(G11), .Z(G1334) );
  HDNAN2D1 U253 ( .A1(n266), .A2(n224), .Z(n267) );
  HDEXOR2D1 U254 ( .A1(n268), .A2(G10), .Z(G1333) );
  HDNAN2D1 U255 ( .A1(n266), .A2(n222), .Z(n268) );
  HDEXOR2D1 U256 ( .A1(n269), .A2(G9), .Z(G1332) );
  HDNAN2D1 U257 ( .A1(n266), .A2(n226), .Z(n269) );
  HDNOR4M1DL U258 ( .A1(n251), .A2(n229), .A3(n235), .A4(n264), .Z(n266) );
  HDNOR2D1 U259 ( .A1(n216), .A2(n218), .Z(n251) );
  HDINVBD1 U260 ( .A(n233), .Z(n218) );
  HDINVBD1 U261 ( .A(n231), .Z(n216) );
  HDEXOR2D1 U262 ( .A1(n270), .A2(G8), .Z(G1331) );
  HDNAN2D1 U263 ( .A1(n271), .A2(n221), .Z(n270) );
  HDEXOR2D1 U264 ( .A1(n272), .A2(G7), .Z(G1330) );
  HDNAN2D1 U265 ( .A1(n271), .A2(n224), .Z(n272) );
  HDEXOR2D1 U266 ( .A1(n273), .A2(G6), .Z(G1329) );
  HDNAN2D1 U267 ( .A1(n271), .A2(n222), .Z(n273) );
  HDEXOR2D1 U268 ( .A1(n274), .A2(G5), .Z(G1328) );
  HDNAN2D1 U269 ( .A1(n271), .A2(n226), .Z(n274) );
  HDNOR4M1DL U270 ( .A1(n250), .A2(n233), .A3(n231), .A4(n264), .Z(n271) );
  HDNOR2D1 U271 ( .A1(n220), .A2(n212), .Z(n250) );
  HDINVBD1 U272 ( .A(n229), .Z(n212) );
  HDINVBD1 U273 ( .A(n235), .Z(n220) );
  HDEXNOR2D1 U274 ( .A1(G4), .A2(n275), .Z(G1327) );
  HDNOR2D1 U275 ( .A1(n253), .A2(n276), .Z(n275) );
  HDEXNOR2D1 U276 ( .A1(G3), .A2(n277), .Z(G1326) );
  HDNOR2D1 U277 ( .A1(n257), .A2(n276), .Z(n277) );
  HDEXNOR2D1 U278 ( .A1(G2), .A2(n278), .Z(G1325) );
  HDNOR2D1 U279 ( .A1(n259), .A2(n276), .Z(n278) );
  HDEXNOR2D1 U280 ( .A1(G1), .A2(n279), .Z(G1324) );
  HDNOR2D1 U281 ( .A1(n262), .A2(n276), .Z(n279) );
  HDNAN3D1 U282 ( .A1(n235), .A2(n231), .A3(n280), .Z(n276) );
  HDNOR3DL U283 ( .A1(n229), .A2(n264), .A3(n233), .Z(n280) );
  HDMUXB2D1 U284 ( .A0(n281), .A1(n282), .SL(n283), .Z(n233) );
  HDEXOR3D1 U285 ( .A1(G22), .A2(G18), .A3(n284), .Z(n283) );
  HDEXOR2D1 U286 ( .A1(G30), .A2(G26), .Z(n284) );
  HDNOR2M1DL U287 ( .A1(n285), .A2(n286), .Z(n282) );
  HDNAN2M1D1 U288 ( .A1(n286), .A2(n285), .Z(n281) );
  HDNAN3D1 U289 ( .A1(G41), .A2(n287), .A3(G38), .Z(n285) );
  HDAOI21D1 U290 ( .A1(G41), .A2(G38), .B(n287), .Z(n286) );
  HDEXOR2D1 U291 ( .A1(n288), .A2(n289), .Z(n287) );
  HDOA33D1 U292 ( .A1(n222), .A2(n242), .A3(n224), .B1(n221), .B2(n236), .B3(
        n226), .Z(n264) );
  HDNOR2D1 U293 ( .A1(n257), .A2(n259), .Z(n236) );
  HDINVBD1 U294 ( .A(n222), .Z(n259) );
  HDINVBD1 U295 ( .A(n224), .Z(n257) );
  HDMUXB2D1 U296 ( .A0(n290), .A1(n291), .SL(n292), .Z(n224) );
  HDEXOR3D1 U297 ( .A1(G15), .A2(G11), .A3(n293), .Z(n292) );
  HDEXOR2D1 U298 ( .A1(G7), .A2(G3), .Z(n293) );
  HDNOR2M1DL U299 ( .A1(n294), .A2(n295), .Z(n291) );
  HDNAN2M1D1 U300 ( .A1(n295), .A2(n294), .Z(n290) );
  HDNAN3D1 U301 ( .A1(G41), .A2(n296), .A3(G35), .Z(n294) );
  HDAOI21D1 U302 ( .A1(G41), .A2(G35), .B(n296), .Z(n295) );
  HDEXOR2D1 U303 ( .A1(n297), .A2(n298), .Z(n296) );
  HDNOR2D1 U304 ( .A1(n262), .A2(n253), .Z(n242) );
  HDINVBD1 U305 ( .A(n221), .Z(n253) );
  HDMUXB2D1 U306 ( .A0(n299), .A1(n300), .SL(n301), .Z(n221) );
  HDEXOR3D1 U307 ( .A1(G16), .A2(G12), .A3(n302), .Z(n301) );
  HDEXOR2D1 U308 ( .A1(G8), .A2(G4), .Z(n302) );
  HDNOR2M1DL U309 ( .A1(n303), .A2(n304), .Z(n300) );
  HDNAN2M1D1 U310 ( .A1(n304), .A2(n303), .Z(n299) );
  HDNAN3D1 U311 ( .A1(G41), .A2(n305), .A3(G36), .Z(n303) );
  HDAOI21D1 U312 ( .A1(G41), .A2(G36), .B(n305), .Z(n304) );
  HDEXNOR2D1 U313 ( .A1(n306), .A2(n307), .Z(n305) );
  HDMUXB2D1 U314 ( .A0(n308), .A1(n309), .SL(n310), .Z(n222) );
  HDEXOR3D1 U315 ( .A1(G14), .A2(G10), .A3(n311), .Z(n310) );
  HDEXOR2D1 U316 ( .A1(G6), .A2(G2), .Z(n311) );
  HDNOR2M1DL U317 ( .A1(n312), .A2(n313), .Z(n309) );
  HDNAN2M1D1 U318 ( .A1(n313), .A2(n312), .Z(n308) );
  HDNAN3D1 U319 ( .A1(G41), .A2(n314), .A3(G34), .Z(n312) );
  HDAOI21D1 U320 ( .A1(G41), .A2(G34), .B(n314), .Z(n313) );
  HDEXNOR2D1 U321 ( .A1(n306), .A2(n297), .Z(n314) );
  HDEXNOR3D1 U322 ( .A1(G26), .A2(G25), .A3(n315), .Z(n297) );
  HDEXNOR2D1 U323 ( .A1(G27), .A2(G28), .Z(n315) );
  HDEXOR3D1 U324 ( .A1(G30), .A2(G29), .A3(n316), .Z(n306) );
  HDEXOR2D1 U325 ( .A1(n214), .A2(G32), .Z(n316) );
  HDINVBD1 U326 ( .A(G31), .Z(n214) );
  HDMUXB2D1 U327 ( .A0(n317), .A1(n318), .SL(n319), .Z(n229) );
  HDEXOR3D1 U328 ( .A1(G24), .A2(G20), .A3(n320), .Z(n319) );
  HDEXOR2D1 U329 ( .A1(G32), .A2(G28), .Z(n320) );
  HDNOR2M1DL U330 ( .A1(n321), .A2(n322), .Z(n318) );
  HDNAN2M1D1 U331 ( .A1(n322), .A2(n321), .Z(n317) );
  HDNAN3D1 U332 ( .A1(G41), .A2(n323), .A3(G40), .Z(n321) );
  HDAOI21D1 U333 ( .A1(G41), .A2(G40), .B(n323), .Z(n322) );
  HDEXOR2D1 U334 ( .A1(n289), .A2(n324), .Z(n323) );
  HDEXOR3D1 U335 ( .A1(G14), .A2(n260), .A3(n325), .Z(n289) );
  HDEXOR2D1 U336 ( .A1(n255), .A2(G16), .Z(n325) );
  HDINVBD1 U337 ( .A(G15), .Z(n255) );
  HDINVBD1 U338 ( .A(G13), .Z(n260) );
  HDMUXB2D1 U339 ( .A0(n326), .A1(n327), .SL(n328), .Z(n231) );
  HDEXOR3D1 U340 ( .A1(G23), .A2(G19), .A3(n329), .Z(n328) );
  HDEXOR2D1 U341 ( .A1(G31), .A2(G27), .Z(n329) );
  HDNOR2M1DL U342 ( .A1(n330), .A2(n331), .Z(n327) );
  HDNAN2M1D1 U343 ( .A1(n331), .A2(n330), .Z(n326) );
  HDNAN3D1 U344 ( .A1(G39), .A2(n332), .A3(G41), .Z(n330) );
  HDAOI21D1 U345 ( .A1(G39), .A2(G41), .B(n332), .Z(n331) );
  HDEXNOR2D1 U346 ( .A1(n333), .A2(n288), .Z(n332) );
  HDEXNOR3D1 U347 ( .A1(G11), .A2(G10), .A3(n334), .Z(n288) );
  HDEXNOR2D1 U348 ( .A1(G12), .A2(G9), .Z(n334) );
  HDMUXB2D1 U349 ( .A0(n335), .A1(n336), .SL(n337), .Z(n235) );
  HDEXOR3D1 U350 ( .A1(G21), .A2(G17), .A3(n338), .Z(n337) );
  HDEXOR2D1 U351 ( .A1(G29), .A2(G25), .Z(n338) );
  HDNOR2M1DL U352 ( .A1(n339), .A2(n340), .Z(n336) );
  HDNAN2M1D1 U353 ( .A1(n340), .A2(n339), .Z(n335) );
  HDNAN3D1 U354 ( .A1(G41), .A2(n341), .A3(G37), .Z(n339) );
  HDAOI21D1 U355 ( .A1(G41), .A2(G37), .B(n341), .Z(n340) );
  HDEXNOR2D1 U356 ( .A1(n333), .A2(n324), .Z(n341) );
  HDEXNOR3D1 U357 ( .A1(G6), .A2(G5), .A3(n342), .Z(n324) );
  HDEXNOR2D1 U358 ( .A1(G7), .A2(G8), .Z(n342) );
  HDEXOR3D1 U359 ( .A1(G2), .A2(G1), .A3(n343), .Z(n333) );
  HDEXNOR2D1 U360 ( .A1(G3), .A2(G4), .Z(n343) );
  HDINVBD1 U361 ( .A(n226), .Z(n262) );
  HDMUXB2D1 U362 ( .A0(n344), .A1(n345), .SL(n346), .Z(n226) );
  HDEXOR3D1 U363 ( .A1(G13), .A2(G1), .A3(n347), .Z(n346) );
  HDEXOR2D1 U364 ( .A1(G9), .A2(G5), .Z(n347) );
  HDNOR2M1DL U365 ( .A1(n348), .A2(n349), .Z(n345) );
  HDNAN2M1D1 U366 ( .A1(n349), .A2(n348), .Z(n344) );
  HDNAN3D1 U367 ( .A1(G41), .A2(n350), .A3(G33), .Z(n348) );
  HDAOI21D1 U368 ( .A1(G41), .A2(G33), .B(n350), .Z(n349) );
  HDEXOR2D1 U369 ( .A1(n298), .A2(n307), .Z(n350) );
  HDEXNOR3D1 U370 ( .A1(G22), .A2(G21), .A3(n351), .Z(n307) );
  HDEXNOR2D1 U371 ( .A1(G23), .A2(G24), .Z(n351) );
  HDEXNOR3D1 U372 ( .A1(G18), .A2(G17), .A3(n352), .Z(n298) );
  HDEXOR2D1 U373 ( .A1(n245), .A2(G20), .Z(n352) );
  HDINVBD1 U374 ( .A(G19), .Z(n245) );
endmodule

