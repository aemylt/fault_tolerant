
module c880 ( N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, 
        N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, 
        N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, 
        N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, 
        N228, N237, N246, N255, N259, N260, N261, N267, N268, N388, N389, N390, 
        N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, 
        N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880 );
  input N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73,
         N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106,
         N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152,
         N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207,
         N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268;
  output N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446,
         N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866,
         N874, N878, N879, N880;
  wire   N276, N290, N291, N292, N297, N342, N344, N351, N353, N354, N356,
         N392, N401, N402, N403, N660, N661, N811, N837, N838, N839, N854,
         N858, N867, N868, N869, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315;
  assign N447 = N276;
  assign N388 = N290;
  assign N389 = N291;
  assign N390 = N292;
  assign N391 = N297;
  assign N418 = N342;
  assign N419 = N344;
  assign N420 = N351;
  assign N421 = N353;
  assign N422 = N354;
  assign N423 = N356;
  assign N446 = N392;
  assign N448 = N401;
  assign N449 = N402;
  assign N450 = N403;
  assign N767 = N660;
  assign N768 = N661;
  assign N850 = N811;
  assign N863 = N837;
  assign N864 = N838;
  assign N865 = N839;
  assign N874 = N854;
  assign N866 = N858;
  assign N878 = N867;
  assign N879 = N868;
  assign N880 = N869;

  HDOAI211DL U167 ( .A1(n178), .A2(n179), .B(n180), .C(n181), .Z(N869) );
  HDAOI222D1 U168 ( .A1(N171), .A2(n182), .B1(N219), .B2(n183), .C1(n184), 
        .C2(N246), .Z(n181) );
  HDOA21DL U169 ( .A1(n185), .A2(n186), .B(n187), .Z(n183) );
  HDOAI211DL U170 ( .A1(n188), .A2(n185), .B(n189), .C(n190), .Z(n187) );
  HDAO21DL U171 ( .A1(n191), .A2(n192), .B(n193), .Z(n189) );
  HDMUXB2D1 U172 ( .A0(N237), .A1(n194), .SL(n195), .Z(n180) );
  HDNOR2D1 U173 ( .A1(n188), .A2(n196), .Z(n194) );
  HDOAI211DL U174 ( .A1(n178), .A2(n197), .B(n198), .C(n199), .Z(N868) );
  HDAOI222D1 U175 ( .A1(N165), .A2(n182), .B1(n200), .B2(N219), .C1(N246), 
        .C2(n201), .Z(n199) );
  HDEXNOR2D1 U176 ( .A1(n202), .A2(n203), .Z(n200) );
  HDNOR2M1DL U177 ( .A1(n204), .A2(n205), .Z(n203) );
  HDMUXB2D1 U178 ( .A0(N237), .A1(n206), .SL(n204), .Z(n198) );
  HDNOR2D1 U179 ( .A1(n205), .A2(n196), .Z(n206) );
  HDINVBD1 U180 ( .A(N91), .Z(n197) );
  HDINVBD1 U181 ( .A(N210), .Z(n178) );
  HDAO211DL U182 ( .A1(n207), .A2(N228), .B(n208), .C(n209), .Z(N867) );
  HDAO22DL U183 ( .A1(N268), .A2(N210), .B1(n210), .B2(N246), .Z(n209) );
  HDOAI22DL U184 ( .A1(n211), .A2(n212), .B1(n213), .B2(n214), .Z(n208) );
  HDAOI21D1 U185 ( .A1(N237), .A2(n210), .B(n182), .Z(n213) );
  HDEXOR2D1 U186 ( .A1(n215), .A2(n207), .Z(n212) );
  HDAOI21D1 U187 ( .A1(n210), .A2(N159), .B(n216), .Z(n207) );
  HDOAI22M10D1 U188 ( .A1(n210), .A2(n214), .B1(n215), .B2(n216), .Z(N858) );
  HDNOR2D1 U189 ( .A1(n210), .A2(N159), .Z(n216) );
  HDOA21DL U190 ( .A1(n202), .A2(n205), .B(n204), .Z(n215) );
  HDNAN2D1 U191 ( .A1(N165), .A2(n201), .Z(n204) );
  HDNOR2D1 U192 ( .A1(n201), .A2(N165), .Z(n205) );
  HDOAI211DL U193 ( .A1(n217), .A2(n218), .B(n219), .C(n220), .Z(n201) );
  HDAOI22D1 U194 ( .A1(N138), .A2(N51), .B1(N96), .B2(n221), .Z(n220) );
  HDNOR2M1DL U195 ( .A1(n186), .A2(n185), .Z(n202) );
  HDINVBD1 U196 ( .A(n195), .Z(n185) );
  HDNAN2D1 U197 ( .A1(N171), .A2(n184), .Z(n195) );
  HDOA21DL U198 ( .A1(n188), .A2(n190), .B(n222), .Z(n186) );
  HDAO211DL U199 ( .A1(n191), .A2(n192), .B(n193), .C(n188), .Z(n222) );
  HDINVBD1 U200 ( .A(n223), .Z(n192) );
  HDINVBD1 U201 ( .A(N177), .Z(n191) );
  HDNOR2D1 U202 ( .A1(n184), .A2(N171), .Z(n188) );
  HDAO211DL U203 ( .A1(N149), .A2(n224), .B(n225), .C(n226), .Z(n184) );
  HDAO22DL U204 ( .A1(N17), .A2(N138), .B1(n221), .B2(N101), .Z(n226) );
  HDAO211DL U205 ( .A1(N143), .A2(n224), .B(n225), .C(n227), .Z(n210) );
  HDAO22DL U206 ( .A1(N8), .A2(N138), .B1(n221), .B2(N91), .Z(n227) );
  HDINVBD1 U207 ( .A(n219), .Z(n225) );
  HDINVBD1 U208 ( .A(n217), .Z(n224) );
  HDAO211DL U209 ( .A1(n228), .A2(N228), .B(n229), .C(n230), .Z(N854) );
  HDAO222DL U210 ( .A1(N177), .A2(n182), .B1(n223), .B2(N246), .C1(N101), .C2(
        N210), .Z(n230) );
  HDOAI22M10D1 U211 ( .A1(N237), .A2(n190), .B1(n211), .B2(n231), .Z(n229) );
  HDEXOR2D1 U212 ( .A1(n193), .A2(n228), .Z(n231) );
  HDAOI21D1 U213 ( .A1(n232), .A2(n233), .B(n234), .Z(n193) );
  HDOA21DL U214 ( .A1(N177), .A2(n223), .B(n190), .Z(n228) );
  HDNAN2D1 U215 ( .A1(N177), .A2(n223), .Z(n190) );
  HDOAI211DL U216 ( .A1(n217), .A2(n235), .B(n219), .C(n236), .Z(n223) );
  HDAOI22D1 U217 ( .A1(N106), .A2(n221), .B1(N152), .B2(N138), .Z(n236) );
  HDNAN2D1 U218 ( .A1(N17), .A2(n237), .Z(n219) );
  HDNAN2M1D1 U219 ( .A1(n238), .A2(N55), .Z(n217) );
  HDNAN4D1 U220 ( .A1(n239), .A2(n240), .A3(n241), .A4(n242), .Z(N839) );
  HDNAN2D1 U221 ( .A1(n182), .A2(N195), .Z(n242) );
  HDAOI32D1 U222 ( .A1(n243), .A2(n244), .A3(N219), .B1(N246), .B2(n245), .Z(
        n241) );
  HDOAI211DL U223 ( .A1(n246), .A2(n247), .B(n248), .C(n249), .Z(n244) );
  HDINVBD1 U224 ( .A(n250), .Z(n247) );
  HDOAI21DL U225 ( .A1(n251), .A2(n252), .B(n250), .Z(n243) );
  HDMUXB2D1 U226 ( .A0(N237), .A1(n253), .SL(n250), .Z(n240) );
  HDNOR2D1 U227 ( .A1(n246), .A2(n196), .Z(n253) );
  HDAOI22D1 U228 ( .A1(N210), .A2(N116), .B1(N260), .B2(N255), .Z(n239) );
  HDNAN3D1 U229 ( .A1(n254), .A2(n255), .A3(n256), .Z(N838) );
  HDAOI222D1 U230 ( .A1(N259), .A2(N255), .B1(n182), .B2(N189), .C1(N210), 
        .C2(N111), .Z(n256) );
  HDAOI22D1 U231 ( .A1(n257), .A2(N219), .B1(n258), .B2(N228), .Z(n255) );
  HDEXNOR2D1 U232 ( .A1(n258), .A2(n259), .Z(n257) );
  HDNOR2D1 U233 ( .A1(n251), .A2(n260), .Z(n259) );
  HDNOR2D1 U234 ( .A1(n261), .A2(n262), .Z(n258) );
  HDAOI22D1 U235 ( .A1(n261), .A2(N237), .B1(N246), .B2(n263), .Z(n254) );
  HDAO211DL U236 ( .A1(n234), .A2(N237), .B(n264), .C(n265), .Z(N837) );
  HDAO222DL U237 ( .A1(N183), .A2(n182), .B1(n266), .B2(N246), .C1(N106), .C2(
        N210), .Z(n265) );
  HDOAI22DL U238 ( .A1(n196), .A2(n267), .B1(n211), .B2(n268), .Z(n264) );
  HDEXOR2D1 U239 ( .A1(n267), .A2(n232), .Z(n268) );
  HDAO21DL U240 ( .A1(n269), .A2(n251), .B(n270), .Z(n232) );
  HDAO21DL U241 ( .A1(n260), .A2(n269), .B(n261), .Z(n270) );
  HDAND2D1 U242 ( .A1(N189), .A2(n263), .Z(n261) );
  HDNAN2M1D1 U243 ( .A1(n252), .A2(n250), .Z(n260) );
  HDNAN2D1 U244 ( .A1(N195), .A2(n245), .Z(n250) );
  HDNOR2D1 U245 ( .A1(n249), .A2(n246), .Z(n252) );
  HDNOR2D1 U246 ( .A1(n248), .A2(n246), .Z(n251) );
  HDNOR2D1 U247 ( .A1(n245), .A2(N195), .Z(n246) );
  HDOAI21DL U248 ( .A1(n271), .A2(n272), .B(n273), .Z(n245) );
  HDAOI21D1 U249 ( .A1(N121), .A2(n221), .B(n274), .Z(n273) );
  HDINVBD1 U250 ( .A(N149), .Z(n272) );
  HDINVBD1 U251 ( .A(n262), .Z(n269) );
  HDNOR2D1 U252 ( .A1(n263), .A2(N189), .Z(n262) );
  HDOAI21DL U253 ( .A1(n271), .A2(n218), .B(n275), .Z(n263) );
  HDAOI21D1 U254 ( .A1(N116), .A2(n221), .B(n274), .Z(n275) );
  HDINVBD1 U255 ( .A(N146), .Z(n218) );
  HDINVBD1 U256 ( .A(N219), .Z(n211) );
  HDNAN2M1D1 U257 ( .A1(n234), .A2(n233), .Z(n267) );
  HDNAN2D1 U258 ( .A1(n276), .A2(n277), .Z(n233) );
  HDNOR2D1 U259 ( .A1(n277), .A2(n276), .Z(n234) );
  HDINVBD1 U260 ( .A(n266), .Z(n276) );
  HDOAI21DL U261 ( .A1(n271), .A2(n278), .B(n279), .Z(n266) );
  HDAOI21D1 U262 ( .A1(N111), .A2(n221), .B(n274), .Z(n279) );
  HDINVBD1 U263 ( .A(N143), .Z(n278) );
  HDNAN3D1 U264 ( .A1(n280), .A2(n281), .A3(n282), .Z(N811) );
  HDAOI222D1 U265 ( .A1(N246), .A2(n283), .B1(n284), .B2(N219), .C1(n182), 
        .C2(N201), .Z(n282) );
  HDAND3D1 U266 ( .A1(N73), .A2(N72), .A3(n285), .Z(n182) );
  HDNOR3DL U267 ( .A1(n286), .A2(n287), .A3(n288), .Z(n285) );
  HDAOI21D1 U268 ( .A1(n289), .A2(n248), .B(n290), .Z(n284) );
  HDMUXB2D1 U269 ( .A0(N237), .A1(n291), .SL(n248), .Z(n281) );
  HDNAN2D1 U270 ( .A1(N201), .A2(n283), .Z(n248) );
  HDAOI21D1 U271 ( .A1(n196), .A2(n292), .B(n293), .Z(n291) );
  HDNAN2D1 U272 ( .A1(N219), .A2(n249), .Z(n292) );
  HDINVBD1 U273 ( .A(n289), .Z(n249) );
  HDNOR2D1 U274 ( .A1(n290), .A2(n293), .Z(n289) );
  HDNOR2D1 U275 ( .A1(n283), .A2(N201), .Z(n293) );
  HDOAI21DL U276 ( .A1(n271), .A2(n235), .B(n294), .Z(n283) );
  HDAOI21D1 U277 ( .A1(N126), .A2(n221), .B(n274), .Z(n294) );
  HDAND2D1 U278 ( .A1(N55), .A2(n237), .Z(n274) );
  HDAND3D1 U279 ( .A1(N80), .A2(N75), .A3(n295), .Z(n237) );
  HDNOR3DL U280 ( .A1(n296), .A2(N268), .A3(n297), .Z(n295) );
  HDOAI21DL U281 ( .A1(n298), .A2(n299), .B(n300), .Z(n221) );
  HDNAN4D1 U282 ( .A1(N59), .A2(N156), .A3(N276), .A4(n301), .Z(n300) );
  HDEXNOR2D1 U283 ( .A1(n288), .A2(N17), .Z(n301) );
  HDOAI31DL U284 ( .A1(n288), .A2(n302), .A3(n287), .B(N51), .Z(n299) );
  HDINVBD1 U285 ( .A(N153), .Z(n235) );
  HDOA21M10D1 U286 ( .A2(n238), .A1(N17), .B(N1), .Z(n271) );
  HDAO21DL U287 ( .A1(N156), .A2(N59), .B(n297), .Z(n238) );
  HDINVBD1 U288 ( .A(N261), .Z(n290) );
  HDINVBD1 U289 ( .A(N228), .Z(n196) );
  HDAOI22D1 U290 ( .A1(N210), .A2(N121), .B1(N267), .B2(N255), .Z(n280) );
  HDEXOR3D1 U291 ( .A1(n303), .A2(n304), .A3(n305), .Z(N661) );
  HDEXOR2D1 U292 ( .A1(N207), .A2(N201), .Z(n305) );
  HDEXNOR3D1 U293 ( .A1(n214), .A2(N130), .A3(n306), .Z(n304) );
  HDEXOR2D1 U294 ( .A1(N171), .A2(N165), .Z(n306) );
  HDINVBD1 U295 ( .A(N159), .Z(n214) );
  HDEXNOR3D1 U296 ( .A1(n277), .A2(N177), .A3(n307), .Z(n303) );
  HDEXOR2D1 U297 ( .A1(N195), .A2(N189), .Z(n307) );
  HDINVBD1 U298 ( .A(N183), .Z(n277) );
  HDEXOR3D1 U299 ( .A1(n308), .A2(n309), .A3(n310), .Z(N660) );
  HDEXOR2D1 U300 ( .A1(N135), .A2(N126), .Z(n310) );
  HDEXOR3D1 U301 ( .A1(N106), .A2(N101), .A3(n311), .Z(n309) );
  HDEXOR2D1 U302 ( .A1(N116), .A2(N111), .Z(n311) );
  HDEXOR3D1 U303 ( .A1(N130), .A2(N121), .A3(n312), .Z(n308) );
  HDEXNOR2D1 U304 ( .A1(n179), .A2(N91), .Z(n312) );
  HDINVBD1 U305 ( .A(N96), .Z(n179) );
  HDNOR2M1DL U306 ( .A1(N89), .A2(n313), .Z(N403) );
  HDNOR3M1DL U307 ( .A1(N74), .A2(n286), .A3(n287), .Z(N402) );
  HDINVBD1 U308 ( .A(N59), .Z(n287) );
  HDNOR2D1 U309 ( .A1(n296), .A2(n286), .Z(N401) );
  HDNAN3D1 U310 ( .A1(N68), .A2(N13), .A3(n314), .Z(n286) );
  HDAND3D1 U311 ( .A1(N8), .A2(N1), .A3(N55), .Z(n314) );
  HDNAN2D1 U312 ( .A1(N292), .A2(n315), .Z(N392) );
  HDNOR2M1DL U313 ( .A1(N90), .A2(n313), .Z(N356) );
  HDNOR2D1 U314 ( .A1(N87), .A2(N88), .Z(n313) );
  HDNAN3D1 U315 ( .A1(N42), .A2(N59), .A3(N36), .Z(N354) );
  HDNAN3D1 U316 ( .A1(N59), .A2(N80), .A3(N36), .Z(N353) );
  HDNAN3D1 U317 ( .A1(N80), .A2(N75), .A3(N59), .Z(N351) );
  HDNAN2M1D1 U318 ( .A1(N292), .A2(n315), .Z(N344) );
  HDAND4D1 U319 ( .A1(N13), .A2(N17), .A3(N26), .A4(N1), .Z(n315) );
  HDNOR2M1DL U320 ( .A1(N13), .A2(n298), .Z(N342) );
  HDNAN3D1 U321 ( .A1(N17), .A2(N1), .A3(N8), .Z(n298) );
  HDAND2D1 U322 ( .A1(N86), .A2(N85), .Z(N297) );
  HDNOR3M1DL U323 ( .A1(N36), .A2(n288), .A3(n296), .Z(N292) );
  HDAND3D1 U324 ( .A1(N36), .A2(N29), .A3(N80), .Z(N291) );
  HDNOR3DL U325 ( .A1(n288), .A2(n296), .A3(n302), .Z(N290) );
  HDINVBD1 U326 ( .A(N75), .Z(n302) );
  HDINVBD1 U327 ( .A(N29), .Z(n296) );
  HDINVBD1 U328 ( .A(N42), .Z(n288) );
  HDINVBD1 U329 ( .A(n297), .Z(N276) );
  HDNAN3D1 U330 ( .A1(N26), .A2(N1), .A3(N51), .Z(n297) );
endmodule

