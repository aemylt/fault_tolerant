
module dff_test_1 ( CK, Q, D, test_si, test_se );
  input CK, D, test_si, test_se;
  output Q;


  HDSDFPQ1 Q_reg ( .D(D), .SD(test_si), .SE(test_se), .CK(CK), .Q(Q) );
endmodule


module dff_test_2 ( CK, Q, D, test_si, test_se );
  input CK, D, test_si, test_se;
  output Q;


  HDSDFPQ1 Q_reg ( .D(D), .SD(test_si), .SE(test_se), .CK(CK), .Q(Q) );
endmodule


module dff_test_3 ( CK, Q, D, test_si, test_se );
  input CK, D, test_si, test_se;
  output Q;


  HDSDFPQ1 Q_reg ( .D(D), .SD(test_si), .SE(test_se), .CK(CK), .Q(Q) );
endmodule


module dff_test_4 ( CK, Q, D, test_si, test_se );
  input CK, D, test_si, test_se;
  output Q;


  HDSDFPQ1 Q_reg ( .D(D), .SD(test_si), .SE(test_se), .CK(CK), .Q(Q) );
endmodule


module dff_test_5 ( CK, Q, D, test_si, test_se );
  input CK, D, test_si, test_se;
  output Q;


  HDSDFPQ1 Q_reg ( .D(D), .SD(test_si), .SE(test_se), .CK(CK), .Q(Q) );
endmodule


module dff_test_6 ( CK, Q, D, test_si, test_se );
  input CK, D, test_si, test_se;
  output Q;


  HDSDFPQ1 Q_reg ( .D(D), .SD(test_si), .SE(test_se), .CK(CK), .Q(Q) );
endmodule


module dff_test_7 ( CK, Q, D, test_si, test_se );
  input CK, D, test_si, test_se;
  output Q;


  HDSDFPQ1 Q_reg ( .D(D), .SD(test_si), .SE(test_se), .CK(CK), .Q(Q) );
endmodule


module dff_test_8 ( CK, Q, D, test_si, test_se );
  input CK, D, test_si, test_se;
  output Q;


  HDSDFPQ1 Q_reg ( .D(D), .SD(test_si), .SE(test_se), .CK(CK), .Q(Q) );
endmodule


module dff_test_9 ( CK, Q, D, test_si, test_se );
  input CK, D, test_si, test_se;
  output Q;


  HDSDFPQ1 Q_reg ( .D(D), .SD(test_si), .SE(test_se), .CK(CK), .Q(Q) );
endmodule


module dff_test_10 ( CK, Q, D, test_si, test_se );
  input CK, D, test_si, test_se;
  output Q;


  HDSDFPQ1 Q_reg ( .D(D), .SD(test_si), .SE(test_se), .CK(CK), .Q(Q) );
endmodule


module dff_test_11 ( CK, Q, D, test_si, test_se );
  input CK, D, test_si, test_se;
  output Q;


  HDSDFPQ1 Q_reg ( .D(D), .SD(test_si), .SE(test_se), .CK(CK), .Q(Q) );
endmodule


module dff_test_12 ( CK, Q, D, test_si, test_se );
  input CK, D, test_si, test_se;
  output Q;


  HDSDFPQ1 Q_reg ( .D(D), .SD(test_si), .SE(test_se), .CK(CK), .Q(Q) );
endmodule


module dff_test_13 ( CK, Q, D, test_si, test_se );
  input CK, D, test_si, test_se;
  output Q;


  HDSDFPQ1 Q_reg ( .D(D), .SD(test_si), .SE(test_se), .CK(CK), .Q(Q) );
endmodule


module dff_test_14 ( CK, Q, D, test_si, test_se );
  input CK, D, test_si, test_se;
  output Q;


  HDSDFPQ1 Q_reg ( .D(D), .SD(test_si), .SE(test_se), .CK(CK), .Q(Q) );
endmodule


module dff_test_15 ( CK, Q, D, test_si, test_se );
  input CK, D, test_si, test_se;
  output Q;


  HDSDFPQ1 Q_reg ( .D(D), .SD(test_si), .SE(test_se), .CK(CK), .Q(Q) );
endmodule


module dff_test_16 ( CK, Q, D, test_si, test_se );
  input CK, D, test_si, test_se;
  output Q;


  HDSDFPQ1 Q_reg ( .D(D), .SD(test_si), .SE(test_se), .CK(CK), .Q(Q) );
endmodule


module dff_test_17 ( CK, Q, D, test_si, test_se );
  input CK, D, test_si, test_se;
  output Q;


  HDSDFPQ1 Q_reg ( .D(D), .SD(test_si), .SE(test_se), .CK(CK), .Q(Q) );
endmodule


module dff_test_18 ( CK, Q, D, test_si, test_se );
  input CK, D, test_si, test_se;
  output Q;


  HDSDFPQ1 Q_reg ( .D(D), .SD(test_si), .SE(test_se), .CK(CK), .Q(Q) );
endmodule


module dff_test_19 ( CK, Q, D, test_si, test_se );
  input CK, D, test_si, test_se;
  output Q;


  HDSDFPQ1 Q_reg ( .D(D), .SD(test_si), .SE(test_se), .CK(CK), .Q(Q) );
endmodule


module dff_test_20 ( CK, Q, D, test_si, test_se );
  input CK, D, test_si, test_se;
  output Q;


  HDSDFPQ1 Q_reg ( .D(D), .SD(test_si), .SE(test_se), .CK(CK), .Q(Q) );
endmodule


module dff_test_21 ( CK, Q, D, test_si, test_se );
  input CK, D, test_si, test_se;
  output Q;


  HDSDFPQ1 Q_reg ( .D(D), .SD(test_si), .SE(test_se), .CK(CK), .Q(Q) );
endmodule


module s382 ( GND, VDD, CK, CLR, FM, GRN1, GRN2, RED1, RED2, TEST, YLW1, YLW2, 
        test_si, test_se );
  input GND, VDD, CK, CLR, FM, TEST, test_si, test_se;
  output GRN1, GRN2, RED1, RED2, YLW1, YLW2;
  wire   TESTL, TESTLVIINLATCHVCDAD, FML, FMLVIINLATCHVCDAD, OLATCH_Y2L,
         TCOMB_YA2, OLATCHVUC_6, Y1C, OLATCHVUC_5, R2C, OLATCH_R1L, OLATCH_G2L,
         TCOMB_GA2, OLATCH_G1L, TCOMB_GA1, OLATCH_FEL, C3_Q3, C3_Q3VD, C3_Q2,
         C3_Q2VD, C3_Q1, C3_Q1VD, C3_Q0, C3_Q0VD, UC_16, UC_16VD, UC_17,
         UC_17VD, UC_18, UC_18VD, UC_19, UC_19VD, UC_8, UC_8VD, UC_9, UC_9VD,
         UC_10, UC_10VD, UC_11, UC_11VD, n2, n49, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207;
  assign YLW2 = OLATCH_Y2L;
  assign RED1 = OLATCH_R1L;
  assign GRN2 = OLATCH_G2L;
  assign GRN1 = OLATCH_G1L;

  dff_test_21 DFF_0 ( .CK(CK), .Q(TESTL), .D(TESTLVIINLATCHVCDAD), .test_si(
        test_si), .test_se(test_se) );
  dff_test_1 DFF_1 ( .CK(CK), .Q(FML), .D(FMLVIINLATCHVCDAD), .test_si(TESTL), 
        .test_se(test_se) );
  dff_test_2 DFF_2 ( .CK(CK), .Q(OLATCH_Y2L), .D(TCOMB_YA2), .test_si(FML), 
        .test_se(test_se) );
  dff_test_3 DFF_3 ( .CK(CK), .Q(OLATCHVUC_6), .D(Y1C), .test_si(OLATCH_Y2L), 
        .test_se(test_se) );
  dff_test_4 DFF_4 ( .CK(CK), .Q(OLATCHVUC_5), .D(R2C), .test_si(OLATCHVUC_6), 
        .test_se(test_se) );
  dff_test_5 DFF_5 ( .CK(CK), .Q(OLATCH_R1L), .D(n49), .test_si(OLATCHVUC_5), 
        .test_se(test_se) );
  dff_test_6 DFF_6 ( .CK(CK), .Q(OLATCH_G2L), .D(TCOMB_GA2), .test_si(
        OLATCH_R1L), .test_se(test_se) );
  dff_test_20 DFF_7 ( .CK(CK), .Q(OLATCH_G1L), .D(TCOMB_GA1), .test_si(UC_11), 
        .test_se(test_se) );
  dff_test_7 DFF_8 ( .CK(CK), .Q(OLATCH_FEL), .D(n2), .test_si(OLATCH_G2L), 
        .test_se(test_se) );
  dff_test_8 DFF_9 ( .CK(CK), .Q(C3_Q3), .D(C3_Q3VD), .test_si(OLATCH_FEL), 
        .test_se(test_se) );
  dff_test_9 DFF_10 ( .CK(CK), .Q(C3_Q2), .D(C3_Q2VD), .test_si(C3_Q3), 
        .test_se(test_se) );
  dff_test_10 DFF_11 ( .CK(CK), .Q(C3_Q1), .D(C3_Q1VD), .test_si(C3_Q2), 
        .test_se(test_se) );
  dff_test_11 DFF_12 ( .CK(CK), .Q(C3_Q0), .D(C3_Q0VD), .test_si(C3_Q1), 
        .test_se(test_se) );
  dff_test_12 DFF_13 ( .CK(CK), .Q(UC_16), .D(UC_16VD), .test_si(C3_Q0), 
        .test_se(test_se) );
  dff_test_13 DFF_14 ( .CK(CK), .Q(UC_17), .D(UC_17VD), .test_si(UC_16), 
        .test_se(test_se) );
  dff_test_14 DFF_15 ( .CK(CK), .Q(UC_18), .D(UC_18VD), .test_si(UC_17), 
        .test_se(test_se) );
  dff_test_15 DFF_16 ( .CK(CK), .Q(UC_19), .D(UC_19VD), .test_si(UC_18), 
        .test_se(test_se) );
  dff_test_16 DFF_17 ( .CK(CK), .Q(UC_8), .D(UC_8VD), .test_si(UC_19), 
        .test_se(test_se) );
  dff_test_17 DFF_18 ( .CK(CK), .Q(UC_9), .D(UC_9VD), .test_si(UC_8), 
        .test_se(test_se) );
  dff_test_18 DFF_19 ( .CK(CK), .Q(UC_10), .D(UC_10VD), .test_si(UC_9), 
        .test_se(test_se) );
  dff_test_19 DFF_20 ( .CK(CK), .Q(UC_11), .D(UC_11VD), .test_si(UC_10), 
        .test_se(test_se) );
  HDOAI31DL U142 ( .A1(n155), .A2(OLATCH_FEL), .A3(C3_Q2), .B(n156), .Z(n49)
         );
  HDAOI21D1 U143 ( .A1(C3_Q0), .A2(n157), .B(n158), .Z(n155) );
  HDINVBD1 U144 ( .A(OLATCHVUC_6), .Z(YLW1) );
  HDOAI21DL U145 ( .A1(n159), .A2(n160), .B(n161), .Z(Y1C) );
  HDOAI31DL U146 ( .A1(n162), .A2(C3_Q1), .A3(C3_Q0), .B(n163), .Z(n161) );
  HDMUXB2D1 U147 ( .A0(n164), .A1(n165), .SL(n158), .Z(n162) );
  HDNOR2D1 U148 ( .A1(n166), .A2(n167), .Z(n165) );
  HDNOR2D1 U149 ( .A1(C3_Q2), .A2(CLR), .Z(n164) );
  HDINVBD1 U150 ( .A(n2), .Z(n159) );
  HDAOI21D1 U151 ( .A1(n168), .A2(n169), .B(n170), .Z(UC_9VD) );
  HDAOI21D1 U152 ( .A1(UC_11), .A2(UC_10), .B(UC_9), .Z(n170) );
  HDNAN2D1 U153 ( .A1(n171), .A2(n172), .Z(n169) );
  HDNOR2D1 U154 ( .A1(n173), .A2(n174), .Z(UC_8VD) );
  HDAOI21D1 U155 ( .A1(n175), .A2(UC_11), .B(UC_8), .Z(n173) );
  HDINVBD1 U156 ( .A(n172), .Z(n175) );
  HDNAN2D1 U157 ( .A1(UC_9), .A2(UC_10), .Z(n172) );
  HDNOR2D1 U158 ( .A1(n176), .A2(n177), .Z(UC_19VD) );
  HDEXNOR2D1 U159 ( .A1(UC_19), .A2(n178), .Z(n177) );
  HDNOR3M1DL U160 ( .A1(n179), .A2(n176), .A3(n180), .Z(UC_18VD) );
  HDAOI21D1 U161 ( .A1(UC_19), .A2(n178), .B(UC_18), .Z(n180) );
  HDAOI211D1 U162 ( .A1(n160), .A2(n179), .B(n176), .C(n181), .Z(UC_17VD) );
  HDAOI21M20D1 U163 ( .A1(UC_16), .A2(n181), .B(n176), .Z(UC_16VD) );
  HDNOR2D1 U164 ( .A1(n179), .A2(n160), .Z(n181) );
  HDNAN3D1 U165 ( .A1(UC_19), .A2(n178), .A3(UC_18), .Z(n179) );
  HDMUXB2D1 U166 ( .A0(n182), .A1(n168), .SL(UC_10), .Z(UC_10VD) );
  HDINVBD1 U167 ( .A(UC_11VD), .Z(n168) );
  HDNOR2D1 U168 ( .A1(n174), .A2(UC_11), .Z(UC_11VD) );
  HDNAN2D1 U169 ( .A1(n171), .A2(UC_11), .Z(n182) );
  HDINVBD1 U170 ( .A(n174), .Z(n171) );
  HDNAN2D1 U171 ( .A1(n183), .A2(n156), .Z(n174) );
  HDNOR2D1 U172 ( .A1(CLR), .A2(n184), .Z(TESTLVIINLATCHVCDAD) );
  HDEXNOR2D1 U173 ( .A1(TESTL), .A2(TEST), .Z(n184) );
  HDNOR3M1DL U174 ( .A1(n185), .A2(OLATCH_FEL), .A3(C3_Q2), .Z(TCOMB_YA2) );
  HDNOR4D1 U175 ( .A1(n185), .A2(n186), .A3(n187), .A4(n188), .Z(TCOMB_GA2) );
  HDAOI211D1 U176 ( .A1(OLATCH_FEL), .A2(n189), .B(n190), .C(n167), .Z(
        TCOMB_GA1) );
  HDOAI21DL U177 ( .A1(n158), .A2(n166), .B(n191), .Z(n190) );
  HDINVBD1 U178 ( .A(OLATCHVUC_5), .Z(RED2) );
  HDMUXB2D1 U179 ( .A0(n192), .A1(n160), .SL(n2), .Z(R2C) );
  HDOAI21DL U180 ( .A1(n167), .A2(n191), .B(n163), .Z(n2) );
  HDOAI21DL U181 ( .A1(n193), .A2(n189), .B(n188), .Z(n163) );
  HDAND2D1 U182 ( .A1(OLATCH_FEL), .A2(n156), .Z(n188) );
  HDNAN4D1 U183 ( .A1(C3_Q0), .A2(n157), .A3(n158), .A4(n166), .Z(n189) );
  HDINVBD1 U184 ( .A(FML), .Z(n166) );
  HDNAN3D1 U185 ( .A1(n194), .A2(n157), .A3(FML), .Z(n191) );
  HDINVBD1 U186 ( .A(UC_17), .Z(n160) );
  HDAO21DL U187 ( .A1(n157), .A2(n186), .B(n187), .Z(n192) );
  HDNOR3DL U188 ( .A1(C3_Q0), .A2(CLR), .A3(n158), .Z(n186) );
  HDNOR2D1 U189 ( .A1(CLR), .A2(n195), .Z(FMLVIINLATCHVCDAD) );
  HDEXNOR2D1 U190 ( .A1(FML), .A2(FM), .Z(n195) );
  HDOAI32DL U191 ( .A1(n196), .A2(n197), .A3(n167), .B1(n158), .B2(n198), .Z(
        C3_Q3VD) );
  HDINVBD1 U192 ( .A(C3_Q3), .Z(n158) );
  HDINVBD1 U193 ( .A(n187), .Z(n167) );
  HDAOI211D1 U194 ( .A1(n199), .A2(C3_Q2), .B(n200), .C(n197), .Z(C3_Q2VD) );
  HDAOI21D1 U195 ( .A1(n201), .A2(n185), .B(n187), .Z(n200) );
  HDNOR2D1 U196 ( .A1(n193), .A2(CLR), .Z(n187) );
  HDNOR3DL U197 ( .A1(n194), .A2(CLR), .A3(n157), .Z(n185) );
  HDNOR3DL U198 ( .A1(n198), .A2(n199), .A3(n202), .Z(C3_Q1VD) );
  HDAOI21D1 U199 ( .A1(n201), .A2(C3_Q0), .B(C3_Q1), .Z(n202) );
  HDINVBD1 U200 ( .A(n196), .Z(n199) );
  HDNAN3D1 U201 ( .A1(C3_Q1), .A2(C3_Q0), .A3(n201), .Z(n196) );
  HDINVBD1 U202 ( .A(n203), .Z(n198) );
  HDMUXB2D1 U203 ( .A0(n176), .A1(n204), .SL(n194), .Z(C3_Q0VD) );
  HDNAN2D1 U204 ( .A1(n203), .A2(n201), .Z(n204) );
  HDNOR2D1 U205 ( .A1(n197), .A2(CLR), .Z(n203) );
  HDAND3D1 U206 ( .A1(n205), .A2(C3_Q3), .A3(n201), .Z(n197) );
  HDINVBD1 U207 ( .A(n206), .Z(n201) );
  HDNAN3D1 U208 ( .A1(n157), .A2(n193), .A3(n194), .Z(n205) );
  HDINVBD1 U209 ( .A(C3_Q0), .Z(n194) );
  HDINVBD1 U210 ( .A(C3_Q2), .Z(n193) );
  HDINVBD1 U211 ( .A(C3_Q1), .Z(n157) );
  HDNAN2D1 U212 ( .A1(n156), .A2(n206), .Z(n176) );
  HDNAN3M1DL U213 ( .A1(n207), .A2(n178), .A3(UC_16), .Z(n206) );
  HDNAN2M1D1 U214 ( .A1(TESTL), .A2(n183), .Z(n178) );
  HDOAI31DL U215 ( .A1(UC_10), .A2(UC_9), .A3(UC_11), .B(UC_8), .Z(n183) );
  HDNOR3DL U216 ( .A1(UC_18), .A2(UC_19), .A3(UC_17), .Z(n207) );
  HDINVBD1 U217 ( .A(CLR), .Z(n156) );
endmodule

